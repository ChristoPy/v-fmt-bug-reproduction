module example

const my_array = [1, 2, 3, 4, 5, 6, 7, 8, 9, 10]

pub fn print_all(example string) {
	for item in my_array {
		println(item)
	}
}
