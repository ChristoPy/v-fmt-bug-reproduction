module main

import example 

fn main() {
	println('Hello World!')
	example.print_all()
}
